// Color drawing
0: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y + 'd2);
end
1: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
2: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
3: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
4: begin
    next_x = $clog2(WIDTH)'(x - 'd2);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
5: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
6: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
7: begin
    next_x = $clog2(WIDTH)'(x - 'd2);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
8: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
9: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
10: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
11: begin
    next_x = $clog2(WIDTH)'(x - 'd3);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
12: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
13: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
14: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
15: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
16: begin
    next_x = $clog2(WIDTH)'(x - 'd4);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
17: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
18: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
19: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
20: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
21: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
22: begin
    next_x = $clog2(WIDTH)'(x - 'd5);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
23: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
24: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
25: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
26: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
27: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
28: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
29: begin
    next_x = $clog2(WIDTH)'(x - 'd6);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
30: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
31: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
32: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
33: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
34: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
35: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
36: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
37: begin
    next_x = $clog2(WIDTH)'(x - 'd7);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
38: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
39: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
40: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
41: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
42: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
43: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
44: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
45: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
46: begin
    next_x = $clog2(WIDTH)'(x - 'd8);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
47: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
48: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
49: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
50: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
51: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
52: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
53: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
54: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
55: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
56: begin
    next_x = $clog2(WIDTH)'(x - 'd9);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
57: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
58: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
59: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
60: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
61: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
62: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
63: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
64: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
65: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
66: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
67: begin
    next_x = $clog2(WIDTH)'(x - 'd10);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
68: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
69: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
70: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
71: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
72: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
73: begin
    next_x = $clog2(WIDTH)'(x - 'd5);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
74: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
75: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
76: begin
    next_x = $clog2(WIDTH)'(x + 'd2);
    next_y = $clog2(HEIGHT)'(y);
end
77: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
78: begin
    next_x = $clog2(WIDTH)'(x - 'd5);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
79: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
80: begin
    next_x = $clog2(WIDTH)'(x + 'd4);
    next_y = $clog2(HEIGHT)'(y);
end
81: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
82: begin
    next_x = $clog2(WIDTH)'(x - 'd6);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
83: begin
    next_x = $clog2(WIDTH)'(x + 'd5);
    next_y = $clog2(HEIGHT)'(y);
end
84: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
85: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
86: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
87: begin
    next_x = $clog2(WIDTH)'(x - 'd1);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
88: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
end
// Black drawing
89: begin
    next_x = $clog2(WIDTH)'(x - 'd8);
    next_y = $clog2(HEIGHT)'(y - 'd18);
    next_color = COLOR_BLACK;
end
90: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
    next_color = COLOR_BLACK;
end
91: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
    next_color = COLOR_BLACK;
end
92: begin
    next_x = $clog2(WIDTH)'(x - 'd1);
    next_y = $clog2(HEIGHT)'(y + 'd1);
    next_color = COLOR_BLACK;
end
93: begin
    next_x = $clog2(WIDTH)'(x + 'd2);
    next_y = $clog2(HEIGHT)'(y);
    next_color = COLOR_BLACK;
end
94: begin
    next_x = $clog2(WIDTH)'(x - 'd2);
    next_y = $clog2(HEIGHT)'(y + 'd1);
    next_color = COLOR_BLACK;
end
95: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
    next_color = COLOR_BLACK;
end
96: begin
    next_x = $clog2(WIDTH)'(x + 'd4);
    next_y = $clog2(HEIGHT)'(y);
    next_color = COLOR_BLACK;
end
97: begin
    next_x = $clog2(WIDTH)'(x - 'd4);
    next_y = $clog2(HEIGHT)'(y + 'd1);
    next_color = COLOR_BLACK;
end
98: begin
    next_x = $clog2(WIDTH)'(x + 'd5);
    next_y = $clog2(HEIGHT)'(y);
    next_color = COLOR_BLACK;
end
99: begin
    next_x = $clog2(WIDTH)'(x - 'd5);
    next_y = $clog2(HEIGHT)'(y + 'd1);
    next_color = COLOR_BLACK;
end
100: begin
    next_x = $clog2(WIDTH)'(x + 'd6);
    next_y = $clog2(HEIGHT)'(y);
    next_color = COLOR_BLACK;
end
101: begin
    next_x = $clog2(WIDTH)'(x - 'd6);
    next_y = $clog2(HEIGHT)'(y + 'd1);
    next_color = COLOR_BLACK;
end
102: begin
    next_x = $clog2(WIDTH)'(x + 'd7);
    next_y = $clog2(HEIGHT)'(y);
    next_color = COLOR_BLACK;
end
103: begin
    next_x = $clog2(WIDTH)'(x - 'd7);
    next_y = $clog2(HEIGHT)'(y + 'd1);
    next_color = COLOR_BLACK;
end
104: begin
    next_x = $clog2(WIDTH)'(x + 'd8);
    next_y = $clog2(HEIGHT)'(y);
    next_color = COLOR_BLACK;
end
105: begin
    next_x = $clog2(WIDTH)'(x - 'd8);
    next_y = $clog2(HEIGHT)'(y + 'd1);
    next_color = COLOR_BLACK;
end
106: begin
    next_x = $clog2(WIDTH)'(x + 'd9);
    next_y = $clog2(HEIGHT)'(y);
    next_color = COLOR_BLACK;
end
107: begin
    next_x = $clog2(WIDTH)'(x - 'd9);
    next_y = $clog2(HEIGHT)'(y + 'd1);
    next_color = COLOR_BLACK;
end
108: begin
    next_x = $clog2(WIDTH)'(x + 'd10);
    next_y = $clog2(HEIGHT)'(y);
    next_color = COLOR_BLACK;
end
109: begin
    next_x = $clog2(WIDTH)'(x - 'd10);
    next_y = $clog2(HEIGHT)'(y + 'd1);
    next_color = COLOR_BLACK;
end
110: begin
    next_x = $clog2(WIDTH)'(x + 'd11);
    next_y = $clog2(HEIGHT)'(y);
    next_color = COLOR_BLACK;
end
111: begin
    next_x = $clog2(WIDTH)'(x - 'd11);
    next_y = $clog2(HEIGHT)'(y + 'd1);
    next_color = COLOR_BLACK;
end
112: begin
    next_x = $clog2(WIDTH)'(x + 'd12);
    next_y = $clog2(HEIGHT)'(y);
    next_color = COLOR_BLACK;
end
113: begin
    next_x = $clog2(WIDTH)'(x - 'd12);
    next_y = $clog2(HEIGHT)'(y + 'd1);
    next_color = COLOR_BLACK;
end
114: begin
    next_x = $clog2(WIDTH)'(x + 'd7);
    next_y = $clog2(HEIGHT)'(y);
    next_color = COLOR_BLACK;
end
115: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
    next_color = COLOR_BLACK;
end
116: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
    next_color = COLOR_BLACK;
end
117: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
    next_color = COLOR_BLACK;
end
118: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
    next_color = COLOR_BLACK;
end
119: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
    next_color = COLOR_BLACK;
end
120: begin
    next_x = $clog2(WIDTH)'(x - 'd12);
    next_y = $clog2(HEIGHT)'(y + 'd1);
    next_color = COLOR_BLACK;
end
121: begin
    next_x = $clog2(WIDTH)'(x + 'd4);
    next_y = $clog2(HEIGHT)'(y);
    next_color = COLOR_BLACK;
end
122: begin
    next_x = $clog2(WIDTH)'(x + 'd3);
    next_y = $clog2(HEIGHT)'(y);
    next_color = COLOR_BLACK;
end
123: begin
    next_x = $clog2(WIDTH)'(x - 'd7);
    next_y = $clog2(HEIGHT)'(y + 'd1);
    next_color = COLOR_BLACK;
end
124: begin
    next_x = $clog2(WIDTH)'(x + 'd3);
    next_y = $clog2(HEIGHT)'(y);
    next_color = COLOR_BLACK;
end
125: begin
    next_x = $clog2(WIDTH)'(x + 'd2);
    next_y = $clog2(HEIGHT)'(y);
    next_color = COLOR_BLACK;
end
126: begin
    next_x = $clog2(WIDTH)'(x + 'd3);
    next_y = $clog2(HEIGHT)'(y);
    next_color = COLOR_BLACK;
end
127: begin
    next_x = $clog2(WIDTH)'(x - 'd8);
    next_y = $clog2(HEIGHT)'(y + 'd1);
    next_color = COLOR_BLACK;
end
128: begin
    next_x = $clog2(WIDTH)'(x + 'd2);
    next_y = $clog2(HEIGHT)'(y);
    next_color = COLOR_BLACK;
end
129: begin
    next_x = $clog2(WIDTH)'(x + 'd3);
    next_y = $clog2(HEIGHT)'(y);
    next_color = COLOR_BLACK;
end
130: begin
    next_x = $clog2(WIDTH)'(x + 'd3);
    next_y = $clog2(HEIGHT)'(y);
    next_color = COLOR_BLACK;
end
131: begin
    next_x = $clog2(WIDTH)'(x - 'd8);
    next_y = $clog2(HEIGHT)'(y + 'd1);
    next_color = COLOR_BLACK;
end
132: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
    next_color = COLOR_BLACK;
end
133: begin
    next_x = $clog2(WIDTH)'(x + 'd5);
    next_y = $clog2(HEIGHT)'(y);
    next_color = COLOR_BLACK;
end
134: begin
    next_x = $clog2(WIDTH)'(x + 'd3);
    next_y = $clog2(HEIGHT)'(y);
    next_color = COLOR_BLACK;
end
135: begin
    next_x = $clog2(WIDTH)'(x - 'd3);
    next_y = $clog2(HEIGHT)'(y + 'd1);
    next_color = COLOR_BLACK;
end
136: begin
    next_x = $clog2(WIDTH)'(x + 'd3);
    next_y = $clog2(HEIGHT)'(y);
    next_color = COLOR_BLACK;
end
137: begin
    next_x = $clog2(WIDTH)'(x - 'd2);
    next_y = $clog2(HEIGHT)'(y + 'd1);
    next_color = COLOR_BLACK;
end
138: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y);
    next_color = COLOR_BLACK;
end
139: begin
    next_x = $clog2(WIDTH)'(x - 'd8);
    next_y = $clog2(HEIGHT)'(y - 'd19);
    next_color = COLOR_BLACK;
end
140: begin
    next_x = x;
    next_y = y;
    next_step = step;
    if (x != cursor_x || y != cursor_y) begin
        next_step = 0;
        ns = STATE_ERASE;
    end
end
default: begin
    next_x = 'x;
    next_y = 'x;
    next_step = 'x;
    $error("Default of STATE_DRAW reached!");
end
