// Erase
0: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y);
end
1: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
2: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
3: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
4: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
5: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
6: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
7: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
8: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
9: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
10: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
11: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
12: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
13: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
14: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
15: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
16: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
17: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
18: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y - 'd16);
end
19: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
20: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
21: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
22: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
23: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
24: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
25: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
26: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
27: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
28: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
29: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
30: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
31: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
32: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
33: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
34: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
35: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y - 'd15);
end
36: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
37: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
38: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
39: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
40: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
41: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
42: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
43: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
44: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
45: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
46: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
47: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
48: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
49: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
50: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y - 'd13);
end
51: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
52: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
53: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
54: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
55: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
56: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
57: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
58: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
59: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
60: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
61: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
62: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
63: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y - 'd11);
end
64: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
65: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
66: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
67: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
68: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
69: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
70: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
71: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
72: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
73: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
74: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y - 'd9);
end
75: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
76: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
77: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
78: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
79: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
80: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
81: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
82: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
83: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
84: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
85: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
86: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y - 'd10);
end
87: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
88: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
89: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
90: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
91: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
92: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
93: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
94: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
95: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
96: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
97: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
98: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
99: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y - 'd11);
end
100: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
101: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
102: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
103: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
104: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
105: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
106: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
107: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
108: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
109: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
110: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
111: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
112: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y - 'd11);
end
113: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
114: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
115: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
116: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
117: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
118: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd2);
end
119: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
120: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
121: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
122: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
123: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y - 'd10);
end
124: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
125: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
126: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
127: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
128: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd4);
end
129: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
130: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y - 'd8);
end
131: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
132: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
133: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
134: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y - 'd2);
end
135: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
136: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
137: begin
    next_x = $clog2(WIDTH)'(x + 'd1);
    next_y = $clog2(HEIGHT)'(y - 'd1);
end
138: begin
    next_x = $clog2(WIDTH)'(x);
    next_y = $clog2(HEIGHT)'(y + 'd1);
end
139: begin
    next_x = x;
    next_y = y;
    next_step = step;
    ns = STATE_INIT;
end
default: begin
    next_x = 'x;
    next_y = 'x;
    next_step = 'x;
    $error("Default of STATE_ERASE reached!");
    $stop;
end
